
2333333333333333333333333333
